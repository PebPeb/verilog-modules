
module MASTER_AXI (
    input clk,

    output AWVALID
  );

  parameter DATA_WIDTH = 32;

  wire clk;

  reg AWVALID = 0;

  always @(posedge clk) begin
    
  end





endmodule
